
module CPU1 (
	clk_clk,
	reset_reset_n,
	leds_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[1:0]	leds_export;
endmodule
