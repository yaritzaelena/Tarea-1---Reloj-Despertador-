
module reloj (
	clk_clk);	

	input		clk_clk;
endmodule
