// reloj_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module reloj_tb (
	);

	wire    reloj_inst_clk_bfm_clk_clk; // reloj_inst_clk_bfm:clk -> reloj_inst:clk_clk

	reloj reloj_inst (
		.clk_clk (reloj_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) reloj_inst_clk_bfm (
		.clk (reloj_inst_clk_bfm_clk_clk)  // clk.clk
	);

endmodule
